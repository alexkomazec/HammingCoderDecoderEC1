library ieee;
use ieee.std_logic_1164.all;

package ram_pkg is
    function clogb2 (depth: in natural) return integer;
end ram_pkg;

package body ram_pkg is

function clogb2( depth : natural) return integer is
variable temp    : integer := depth;
variable ret_val : integer := 0;
begin
    while temp > 1 loop
        ret_val := ret_val + 1;
        temp    := temp / 2;
    end loop;
    return ret_val;
end function;

end package body ram_pkg;

library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.ram_pkg.all;

entity RAM_14bits is
generic (
    RAM_WIDTH : integer:= 14;                      
    RAM_DEPTH : integer:= 292                      
    );

port (
        addra : in std_logic_vector((clogb2(RAM_DEPTH)-1) downto 0);
        dina  : in std_logic_vector(RAM_WIDTH-1 downto 0);		            
        clka  : in std_logic;                       			            
        wea   : in std_logic;                       			            
        douta : out std_logic_vector(RAM_WIDTH-1 downto 0)   			    
    );

end RAM_14bits;

architecture rtl of RAM_14bits is

constant C_RAM_WIDTH : integer := RAM_WIDTH;
constant C_RAM_DEPTH : integer := RAM_DEPTH;

type ram_type is array (C_RAM_DEPTH-1 downto 0) of std_logic_vector (C_RAM_WIDTH-1 downto 0);          
signal ram_name : ram_type:=
    ("00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000",
     "00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000","00000000000000");

begin

process(clka)
begin
    if(clka'event and clka = '1') then
            if(wea = '1') then
                ram_name(to_integer(unsigned(addra(3 downto 0)))) <= dina;
            else
                douta <= ram_name(to_integer(unsigned(addra(3 downto 0))));
            end if;
    end if;
end process;

end rtl;


						
						